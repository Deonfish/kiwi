module Operands(
	input clk,
	input rst_n,
	// stall from scoreboard
	input stall_operands_i,
	// flush from wb
	input flush_operands_i,
	// from decoder
	input [0:0]  inst0_decoder_valid_i,
	input [63:0] inst0_pc_i,
	input [31:0] inst0_inst_i,
	input [0:0]  inst0_rs1_valid_i,
	input [4:0]  inst0_rs1_i,
	input [0:0]  inst0_rs2_valid_i,
	input [4:0]  inst0_rs2_i,
	input [0:0]  inst0_rs3_valid_i,
	input [4:0]  inst0_rs3_i,
	input [1:0]  inst0_rd_type_i,
	input [4:0]  inst0_rd_i,
	input [5:0]  inst0_exe_unit_i,
	input [3:0]  inst0_func_code_i,
	input [2:0]  inst0_func3_i,
	input [1:0]  inst0_func2_i,
	input [0:0]  inst0_endsim_i,
	input [0:0]  inst0_auipc_i,
	input [0:0]  inst1_decoder_valid_i,
	input [63:0] inst1_pc_i,
	input [31:0] inst1_inst_i,
	input [0:0]  inst1_rs1_valid_i,
	input [4:0]  inst1_rs1_i,
	input [0:0]  inst1_rs2_valid_i,
	input [4:0]  inst1_rs2_i,
	input [0:0]  inst1_rs3_valid_i,
	input [4:0]  inst1_rs3_i,
	input [1:0]  inst1_rd_type_i,
	input [4:0]  inst1_rd_i,
	input [5:0]  inst1_exe_unit_i,
	input [3:0]  inst1_func_code_i,
	input [2:0]  inst1_func3_i,
	input [1:0]  inst1_func2_i,
	input [0:0]  inst1_endsim_i,
	input [0:0]  inst1_auipc_i,
	// to operands
	output [0:0]  inst0_operands_valid_o,
	output [63:0] inst0_pc_o,
	output [31:0] inst0_inst_o,
	output [0:0]  inst0_rs1_valid_o,
	output [4:0]  inst0_rs1_o,
	output [63:0] inst0_rs1_value_o,
	output [0:0]  inst0_rs2_valid_o,
	output [4:0]  inst0_rs2_o,
	output [63:0] inst0_rs2_value_o,
	output [0:0]  inst0_rs3_valid_o,
	output [4:0]  inst0_rs3_o,
	output [63:0] inst0_rs3_value_o,
	output [1:0]  inst0_rd_type_o,
	output [4:0]  inst0_rd_o,
	output [5:0]  inst0_exe_unit_o,
	output [3:0]  inst0_func_code_o,
	output [2:0]  inst0_func3_o,
	output [1:0]  inst0_func2_o,
	output [0:0]  inst0_endsim_o,
	output [0:0]  inst0_auipc_o,
	output [0:0]  inst1_operands_valid_o,
	output [63:0] inst1_pc_o,
	output [31:0] inst1_inst_o,
	output [0:0]  inst1_rs1_valid_o,
	output [4:0]  inst1_rs1_o,
	output [63:0] inst1_rs1_value_o,
	output [0:0]  inst1_rs2_valid_o,
	output [4:0]  inst1_rs2_o,
	output [63:0] inst1_rs2_value_o,
	output [0:0]  inst1_rs3_valid_o,
	output [4:0]  inst1_rs3_o,
	output [63:0] inst1_rs3_value_o,
	output [1:0]  inst1_rd_type_o,
	output [4:0]  inst1_rd_o,
	output [5:0]  inst1_exe_unit_o,
	output [3:0]  inst1_func_code_o,
	output [2:0]  inst1_func3_o,
	output [1:0]  inst1_func2_o,
	output [0:0]  inst1_endsim_o,
	output [0:0]  inst1_auipc_o,
    // write reg from wb
    input [0:0]  inst0_wb_valid_i,
    input [4:0]  inst0_wb_rd_i,
    input [63:0] inst0_wb_value_i,
    input [0:0]  inst1_wb_valid_i,
    input [4:0]  inst1_wb_rd_i,
    input [63:0] inst1_wb_value_i
);

module Regfile (
	input 		  clk,
	input 		  rst_n,
	// read
	input [4:0]   inst0_rs1_addr_i,
	input [4:0]   inst0_rs2_addr_i,
	input [4:0]   inst0_rd_addr_i,
	output [63:0] inst0_rs1_rdata_o,
	output [63:0] inst0_rs2_rdata_o,
	output [63:0] inst0_rd_rdata_o,
	input [4:0]   inst1_rs1_addr_i,
	input [4:0]   inst1_rs2_addr_i,
	input [4:0]   inst1_rd_addr_i,
	output [63:0] inst1_rs1_rdata_o,
	output [63:0] inst1_rs2_rdata_o,
	output [63:0] inst1_rd_rdata_o,
	// write
	input [0:0]  inst0_rd_wvalid_i,
	input [4:0]  inst0_rd_waddr_i,
	input [63:0] inst0_rd_wdata_i,
	input [0:0]  inst1_rd_wvalid_i,
	input [4:0]  inst1_rd_waddr_i,
	input [63:0] inst1_rd_wdata_i
);

Regfile u_regfile(
    .clk(clk),
    .rst_n(rst_n),
    .inst0_rs1_addr_i(inst0_rs1_i),
    .inst0_rs2_addr_i(inst0_rs2_i),
    .inst0_rd_addr_i(inst0_rd_i),
    .inst1_rs1_addr_i(inst1_rs1_i),
    .inst1_rs2_addr_i(inst1_rs2_i),
    .inst1_rd_addr_i(inst1_rd_i),
    .inst0_rd_wvalid_i(inst0_wb_valid_i),
    .inst0_rd_waddr_i(inst0_wb_rd_i),
    .inst0_rd_wdata_i(inst0_wb_value_i),
    .inst1_rd_wvalid_i(inst1_wb_valid_i),
    .inst1_rd_waddr_i(inst1_wb_rd_i),
    .inst1_rd_wdata_i(inst1_wb_value_i)
)

endmodule